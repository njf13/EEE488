* Netlist for Tree
* Netlist created on 10:53:21.326 PM 15-Apr-2019

.param maxV = 10


.op
*Vsource Vsource gnd {maxV} AC 1
*.AC dec 10 10 1G
.tran 1ns 1
Vsource Vsource gnd PULSE (0 {maxV} 0 1n 1n 99m 200m)
.measure tran tdlay TRIG V(Vsource) VAL = 0.5*maxV RISE=3 TARG V(n2) VAL = 0.5*maxV RISE=3

Vgnd n1 gnd 0

r1 n1 n2 6.554545454545454
c1 n2 gnd 793.0999999999999u
r2 n2 n3 5.78075068436666
c2 n3 gnd 440.63842899999986u
r3 n2 n4 5.78075068436666
c3 n4 gnd 440.63842899999986u
r4 n4 n6 5.0983060086388585
c4 n6 gnd 244.8143047681099u
r5 n4 n5 5.0983060086388585
c5 n5 gnd 244.8143047681099u
r6 n3 n8 5.0983060086388585
c6 n8 gnd 244.8143047681099u
r7 n3 n7 5.0983060086388585
c7 n7 gnd 244.8143047681099u
r8 n8 n10 4.4964271211379625
c8 n10 gnd 136.01637958611417u
r9 n8 n9 4.4964271211379625
c9 n9 gnd 136.01637958611417u
r10 n6 n12 4.4964271211379625
c10 n12 gnd 136.01637958611417u
r11 n5 n16 4.4964271211379625
c11 n16 gnd 136.01637958611417u
r12 n7 n14 4.4964271211379625
c12 n14 gnd 136.01637958611417u
r13 n7 n13 4.4964271211379625
c13 n13 gnd 136.01637958611417u
r14 n5 n15 4.4964271211379625
c14 n15 gnd 136.01637958611417u
r15 n6 n11 4.4964271211379625
c15 n11 gnd 136.01637958611417u
r16 n10 n20 3.965602853466767
c16 n20 gnd 75.56934033424916u
r17 n10 n19 3.965602853466767
c17 n19 gnd 75.56934033424916u
r18 n15 n32 3.965602853466767
c18 n32 gnd 75.56934033424916u
r19 n13 n23 3.965602853466767
c19 n23 gnd 75.56934033424916u
r21 n9 n22 3.965602853466767
c21 n22 gnd 75.56934033424916u
r22 n11 n25 3.965602853466767
c22 n25 gnd 75.56934033424916u
r23 n16 n17 3.965602853466767
c23 n17 gnd 75.56934033424916u
r24 n11 n26 3.965602853466767
c24 n26 gnd 75.56934033424916u
r25 n13 n24 3.965602853466767
c25 n24 gnd 75.56934033424916u
r26 n16 n18 3.965602853466767
c26 n18 gnd 75.56934033424916u
r27 n12 n29 3.965602853466767
c27 n29 gnd 75.56934033424916u
r28 n14 n28 3.965602853466767
c28 n28 gnd 75.56934033424916u
r29 n12 n30 3.965602853466767
c29 n30 gnd 75.56934033424916u
r30 n14 n27 3.965602853466767
c30 n27 gnd 75.56934033424916u
r31 n9 n21 3.965602853466767
c31 n21 gnd 75.56934033424916u
r32 n24 n56 3.497444875175428
c32 n56 gnd 41.98556979630549u
r33 n29 n61 3.497444875175428
c33 n61 gnd 41.98556979630549u
r34 n22 n39 3.497444875175428
c34 n39 gnd 41.98556979630549u
r35 n17 n37 3.497444875175428
c35 n37 gnd 41.98556979630549u
r36 n23 n34 3.497444875175428
c36 n34 gnd 41.98556979630549u
r37 n21 n43 3.497444875175428
c37 n43 gnd 41.98556979630549u
r39 n30 n36 3.497444875175428
c39 n36 gnd 41.98556979630549u
r40 n20 n47 3.497444875175428
c40 n47 gnd 41.98556979630549u
r41 n23 n33 3.497444875175428
c41 n33 gnd 41.98556979630549u
r42 n25 n51 3.497444875175428
c42 n51 gnd 41.98556979630549u
r43 n29 n62 3.497444875175428
c43 n62 gnd 41.98556979630549u
r44 n26 n45 3.497444875175428
c44 n45 gnd 41.98556979630549u
r45 n22 n40 3.497444875175428
c45 n40 gnd 41.98556979630549u
r47 n17 n38 3.497444875175428
c47 n38 gnd 41.98556979630549u
r48 n21 n44 3.497444875175428
c48 n44 gnd 41.98556979630549u
r49 n18 n57 3.497444875175428
c49 n57 gnd 41.98556979630549u
r50 n26 n46 3.497444875175428
c50 n46 gnd 41.98556979630549u
r51 n32 n54 3.497444875175428
c51 n54 gnd 41.98556979630549u
r52 n24 n55 3.497444875175428
c52 n55 gnd 41.98556979630549u
r54 n19 n60 3.497444875175428
c54 n60 gnd 41.98556979630549u
r55 n27 n50 3.497444875175428
c55 n50 gnd 41.98556979630549u
r56 n30 n35 3.497444875175428
c56 n35 gnd 41.98556979630549u
r57 n19 n59 3.497444875175428
c57 n59 gnd 41.98556979630549u
r58 n27 n49 3.497444875175428
c58 n49 gnd 41.98556979630549u
r60 n25 n52 3.497444875175428
c60 n52 gnd 41.98556979630549u
r61 n28 n41 3.497444875175428
c61 n41 gnd 41.98556979630549u
r62 n37 n99 3.084555137486203
c62 n99 gnd 23.326762723129363u
r63 n60 n72 3.084555137486203
c63 n72 gnd 23.326762723129363u
r64 n40 n83 3.084555137486203
c64 n83 gnd 23.326762723129363u
r65 n38 n96 3.084555137486203
c65 n96 gnd 23.326762723129363u
r66 n61 n101 3.084555137486203
c66 n101 gnd 23.326762723129363u
r67 n56 n86 3.084555137486203
c67 n86 gnd 23.326762723129363u
r68 n33 n63 3.084555137486203
c68 n63 gnd 23.326762723129363u
r69 n50 n110 3.084555137486203
c69 n110 gnd 23.326762723129363u
r70 n52 n65 3.084555137486203
c70 n65 gnd 23.326762723129363u
r71 n45 n73 3.084555137486203
c71 n73 gnd 23.326762723129363u
r72 n36 n87 3.084555137486203
c72 n87 gnd 23.326762723129363u
r73 n45 n74 3.084555137486203
c73 n74 gnd 23.326762723129363u
r74 n55 n91 3.084555137486203
c74 n91 gnd 23.326762723129363u
r75 n36 n88 3.084555137486203
c75 n88 gnd 23.326762723129363u
r76 n60 n71 3.084555137486203
c76 n71 gnd 23.326762723129363u
r77 n61 n102 3.084555137486203
c77 n102 gnd 23.326762723129363u
r78 n49 n80 3.084555137486203
c78 n80 gnd 23.326762723129363u
r79 n54 n81 3.084555137486203
c79 n81 gnd 23.326762723129363u
r82 n37 n100 3.084555137486203
c82 n100 gnd 23.326762723129363u
r83 n35 n67 3.084555137486203
c83 n67 gnd 23.326762723129363u
r84 n39 n89 3.084555137486203
c84 n89 gnd 23.326762723129363u
r85 n52 n66 3.084555137486203
c85 n66 gnd 23.326762723129363u
r86 n40 n84 3.084555137486203
c86 n84 gnd 23.326762723129363u
r87 n57 n93 3.084555137486203
c87 n93 gnd 23.326762723129363u
r88 n46 n111 3.084555137486203
c88 n111 gnd 23.326762723129363u
r90 n62 n98 3.084555137486203
c90 n98 gnd 23.326762723129363u
r91 n34 n105 3.084555137486203
c91 n105 gnd 23.326762723129363u
r93 n57 n94 3.084555137486203
c93 n94 gnd 23.326762723129363u
r94 n62 n97 3.084555137486203
c94 n97 gnd 23.326762723129363u
r95 n38 n95 3.084555137486203
c95 n95 gnd 23.326762723129363u
r97 n55 n92 3.084555137486203
c97 n92 gnd 23.326762723129363u
r98 n50 n109 3.084555137486203
c98 n109 gnd 23.326762723129363u
r100 n34 n106 3.084555137486203
c100 n106 gnd 23.326762723129363u
r101 n44 n75 3.084555137486203
c101 n75 gnd 23.326762723129363u
r103 n59 n70 3.084555137486203
c103 n70 gnd 23.326762723129363u
r104 n35 n68 3.084555137486203
c104 n68 gnd 23.326762723129363u
r105 n41 n114 3.084555137486203
c105 n114 gnd 23.326762723129363u
r106 n56 n85 3.084555137486203
c106 n85 gnd 23.326762723129363u
r107 n44 n76 3.084555137486203
c107 n76 gnd 23.326762723129363u
r109 n33 n64 3.084555137486203
c109 n64 gnd 23.326762723129363u
r110 n41 n113 3.084555137486203
c110 n113 gnd 23.326762723129363u
r111 n39 n90 3.084555137486203
c111 n90 gnd 23.326762723129363u
r112 n47 n103 3.084555137486203
c112 n103 gnd 23.326762723129363u
r114 n65 n147 2.7204089659069446
c114 n147 gnd 12.960116101343441u
r115 n71 n129 2.7204089659069446
c115 n129 gnd 12.960116101343441u
r116 n103 n137 2.7204089659069446
c116 n137 gnd 12.960116101343441u
r117 n113 n166 2.7204089659069446
c117 n166 gnd 12.960116101343441u
r118 n91 n152 2.7204089659069446
c118 n152 gnd 12.960116101343441u
r119 n70 n174 2.7204089659069446
c119 n174 gnd 12.960116101343441u
r120 n89 n178 2.7204089659069446
c120 n178 gnd 12.960116101343441u
r121 n67 n143 2.7204089659069446
c121 n143 gnd 12.960116101343441u
r122 n73 n131 2.7204089659069446
c122 n131 gnd 12.960116101343441u
r123 n97 n140 2.7204089659069446
c123 n140 gnd 12.960116101343441u
r126 n109 n170 2.7204089659069446
c126 n170 gnd 12.960116101343441u
r128 n70 n173 2.7204089659069446
c128 n173 gnd 12.960116101343441u
r130 n96 n182 2.7204089659069446
c130 n182 gnd 12.960116101343441u
r131 n74 n184 2.7204089659069446
c131 n184 gnd 12.960116101343441u
r132 n114 n161 2.7204089659069446
c132 n161 gnd 12.960116101343441u
r133 n81 n157 2.7204089659069446
c133 n157 gnd 12.960116101343441u
r134 n95 n191 2.7204089659069446
c134 n191 gnd 12.960116101343441u
r135 n92 n128 2.7204089659069446
c135 n128 gnd 12.960116101343441u
r136 n105 n145 2.7204089659069446
c136 n145 gnd 12.960116101343441u
r137 n87 n194 2.7204089659069446
c137 n194 gnd 12.960116101343441u
r138 n74 n183 2.7204089659069446
c138 n183 gnd 12.960116101343441u
r139 n110 n164 2.7204089659069446
c139 n164 gnd 12.960116101343441u
r140 n85 n187 2.7204089659069446
c140 n187 gnd 12.960116101343441u
r141 n63 n200 2.7204089659069446
c141 n200 gnd 12.960116101343441u
r142 n114 n162 2.7204089659069446
c142 n162 gnd 12.960116101343441u
r143 n90 n122 2.7204089659069446
c143 n122 gnd 12.960116101343441u
r145 n73 n132 2.7204089659069446
c145 n132 gnd 12.960116101343441u
r146 n68 n168 2.7204089659069446
c146 n168 gnd 12.960116101343441u
r147 n111 n124 2.7204089659069446
c147 n124 gnd 12.960116101343441u
r151 n71 n130 2.7204089659069446
c151 n130 gnd 12.960116101343441u
r152 n66 n117 2.7204089659069446
c152 n117 gnd 12.960116101343441u
r153 n67 n144 2.7204089659069446
c153 n144 gnd 12.960116101343441u
r154 n76 n195 2.7204089659069446
c154 n195 gnd 12.960116101343441u
r155 n109 n169 2.7204089659069446
c155 n169 gnd 12.960116101343441u
r157 n96 n181 2.7204089659069446
c157 n181 gnd 12.960116101343441u
r159 n75 n186 2.7204089659069446
c159 n186 gnd 12.960116101343441u
r160 n98 n133 2.7204089659069446
c160 n133 gnd 12.960116101343441u
r161 n91 n151 2.7204089659069446
c161 n151 gnd 12.960116101343441u
r162 n88 n135 2.7204089659069446
c162 n135 gnd 12.960116101343441u
r164 n72 n155 2.7204089659069446
c164 n155 gnd 12.960116101343441u
r165 n97 n139 2.7204089659069446
c165 n139 gnd 12.960116101343441u
r167 n81 n158 2.7204089659069446
c167 n158 gnd 12.960116101343441u
r168 n80 n175 2.7204089659069446
c168 n175 gnd 12.960116101343441u
r169 n64 n141 2.7204089659069446
c169 n141 gnd 12.960116101343441u
r170 n80 n176 2.7204089659069446
c170 n176 gnd 12.960116101343441u
r171 n64 n142 2.7204089659069446
c171 n142 gnd 12.960116101343441u
r172 n106 n197 2.7204089659069446
c172 n197 gnd 12.960116101343441u
r173 n87 n193 2.7204089659069446
c173 n193 gnd 12.960116101343441u
r174 n102 n180 2.7204089659069446
c174 n180 gnd 12.960116101343441u
r175 n83 n189 2.7204089659069446
c175 n189 gnd 12.960116101343441u
r176 n63 n199 2.7204089659069446
c176 n199 gnd 12.960116101343441u
r178 n68 n167 2.7204089659069446
c178 n167 gnd 12.960116101343441u
r179 n65 n148 2.7204089659069446
c179 n148 gnd 12.960116101343441u
r181 n105 n146 2.7204089659069446
c181 n146 gnd 12.960116101343441u
r182 n110 n163 2.7204089659069446
c182 n163 gnd 12.960116101343441u
r183 n111 n123 2.7204089659069446
c183 n123 gnd 12.960116101343441u
r185 n88 n136 2.7204089659069446
c185 n136 gnd 12.960116101343441u
r186 n83 n190 2.7204089659069446
c186 n190 gnd 12.960116101343441u
r188 n90 n121 2.7204089659069446
c188 n121 gnd 12.960116101343441u
r189 n103 n138 2.7204089659069446
c189 n138 gnd 12.960116101343441u
r190 n94 n153 2.7204089659069446
c190 n153 gnd 12.960116101343441u
r191 n100 n120 2.7204089659069446
c191 n120 gnd 12.960116101343441u
r192 n92 n127 2.7204089659069446
c192 n127 gnd 12.960116101343441u
r193 n93 n172 2.7204089659069446
c193 n172 gnd 12.960116101343441u
r194 n102 n179 2.7204089659069446
c194 n179 gnd 12.960116101343441u
r196 n95 n192 2.7204089659069446
c196 n192 gnd 12.960116101343441u
r197 n100 n119 2.7204089659069446
c197 n119 gnd 12.960116101343441u
r199 n85 n188 2.7204089659069446
c199 n188 gnd 12.960116101343441u
r200 n124 Vsource 2.399251954308758
c200 Vsource gnd 7.200510904745402u
r201 n168 Vsource 2.399251954308758
c201 Vsource gnd 7.200510904745402u
r202 n153 Vsource 2.399251954308758
c202 Vsource gnd 7.200510904745402u
r203 n191 Vsource 2.399251954308758
c203 Vsource gnd 7.200510904745402u
r204 n127 Vsource 2.399251954308758
c204 Vsource gnd 7.200510904745402u
r205 n197 Vsource 2.399251954308758
c205 Vsource gnd 7.200510904745402u
r206 n200 Vsource 2.399251954308758
c206 Vsource gnd 7.200510904745402u
r207 n181 Vsource 2.399251954308758
c207 Vsource gnd 7.200510904745402u
r208 n184 Vsource 2.399251954308758
c208 Vsource gnd 7.200510904745402u
r209 n183 Vsource 2.399251954308758
c209 Vsource gnd 7.200510904745402u
r210 n129 Vsource 2.399251954308758
c210 Vsource gnd 7.200510904745402u
r211 n187 Vsource 2.399251954308758
c211 Vsource gnd 7.200510904745402u
r212 n180 Vsource 2.399251954308758
c212 Vsource gnd 7.200510904745402u
r213 n178 Vsource 2.399251954308758
c213 Vsource gnd 7.200510904745402u
r214 n170 Vsource 2.399251954308758
c214 Vsource gnd 7.200510904745402u
r215 n131 Vsource 2.399251954308758
c215 Vsource gnd 7.200510904745402u
r216 n190 Vsource 2.399251954308758
c216 Vsource gnd 7.200510904745402u
r217 n190 Vsource 2.399251954308758
c217 Vsource gnd 7.200510904745402u
r218 n121 Vsource 2.399251954308758
c218 Vsource gnd 7.200510904745402u
r220 n191 Vsource 2.399251954308758
c220 Vsource gnd 7.200510904745402u
r221 n199 Vsource 2.399251954308758
c221 Vsource gnd 7.200510904745402u
r222 n162 Vsource 2.399251954308758
c222 Vsource gnd 7.200510904745402u
r223 n170 Vsource 2.399251954308758
c223 Vsource gnd 7.200510904745402u
r224 n167 Vsource 2.399251954308758
c224 Vsource gnd 7.200510904745402u
r226 n135 Vsource 2.399251954308758
c226 Vsource gnd 7.200510904745402u
r227 n141 Vsource 2.399251954308758
c227 Vsource gnd 7.200510904745402u
r229 n130 Vsource 2.399251954308758
c229 Vsource gnd 7.200510904745402u
r230 n128 Vsource 2.399251954308758
c230 Vsource gnd 7.200510904745402u
r231 n169 Vsource 2.399251954308758
c231 Vsource gnd 7.200510904745402u
r232 n167 Vsource 2.399251954308758
c232 Vsource gnd 7.200510904745402u
r233 n161 Vsource 2.399251954308758
c233 Vsource gnd 7.200510904745402u
r234 n189 Vsource 2.399251954308758
c234 Vsource gnd 7.200510904745402u
r235 n164 Vsource 2.399251954308758
c235 Vsource gnd 7.200510904745402u
r236 n155 Vsource 2.399251954308758
c236 Vsource gnd 7.200510904745402u
r237 n145 Vsource 2.399251954308758
c237 Vsource gnd 7.200510904745402u
r238 n145 Vsource 2.399251954308758
c238 Vsource gnd 7.200510904745402u
r239 n184 Vsource 2.399251954308758
c239 Vsource gnd 7.200510904745402u
r240 n195 Vsource 2.399251954308758
c240 Vsource gnd 7.200510904745402u
r241 n135 Vsource 2.399251954308758
c241 Vsource gnd 7.200510904745402u
r242 n163 Vsource 2.399251954308758
c242 Vsource gnd 7.200510904745402u
r243 n192 Vsource 2.399251954308758
c243 Vsource gnd 7.200510904745402u
r244 n148 Vsource 2.399251954308758
c244 Vsource gnd 7.200510904745402u
r246 n148 Vsource 2.399251954308758
c246 Vsource gnd 7.200510904745402u
r248 n140 Vsource 2.399251954308758
c248 Vsource gnd 7.200510904745402u
r249 n166 Vsource 2.399251954308758
c249 Vsource gnd 7.200510904745402u
r250 n127 Vsource 2.399251954308758
c250 Vsource gnd 7.200510904745402u
r251 n197 Vsource 2.399251954308758
c251 Vsource gnd 7.200510904745402u
r253 n124 Vsource 2.399251954308758
c253 Vsource gnd 7.200510904745402u
r254 n152 Vsource 2.399251954308758
c254 Vsource gnd 7.200510904745402u
r255 n123 Vsource 2.399251954308758
c255 Vsource gnd 7.200510904745402u
r256 n132 Vsource 2.399251954308758
c256 Vsource gnd 7.200510904745402u
r259 n119 Vsource 2.399251954308758
c259 Vsource gnd 7.200510904745402u
r260 n133 Vsource 2.399251954308758
c260 Vsource gnd 7.200510904745402u
r261 n192 Vsource 2.399251954308758
c261 Vsource gnd 7.200510904745402u
r264 n174 Vsource 2.399251954308758
c264 Vsource gnd 7.200510904745402u
r265 n195 Vsource 2.399251954308758
c265 Vsource gnd 7.200510904745402u
r266 n193 Vsource 2.399251954308758
c266 Vsource gnd 7.200510904745402u
r267 n136 Vsource 2.399251954308758
c267 Vsource gnd 7.200510904745402u
r268 n121 Vsource 2.399251954308758
c268 Vsource gnd 7.200510904745402u
r269 n176 Vsource 2.399251954308758
c269 Vsource gnd 7.200510904745402u
r270 n194 Vsource 2.399251954308758
c270 Vsource gnd 7.200510904745402u
r272 n182 Vsource 2.399251954308758
c272 Vsource gnd 7.200510904745402u
r273 n178 Vsource 2.399251954308758
c273 Vsource gnd 7.200510904745402u
r275 n189 Vsource 2.399251954308758
c275 Vsource gnd 7.200510904745402u
r276 n183 Vsource 2.399251954308758
c276 Vsource gnd 7.200510904745402u
r277 n136 Vsource 2.399251954308758
c277 Vsource gnd 7.200510904745402u
r280 n186 Vsource 2.399251954308758
c280 Vsource gnd 7.200510904745402u
r283 n158 Vsource 2.399251954308758
c283 Vsource gnd 7.200510904745402u
r284 n163 Vsource 2.399251954308758
c284 Vsource gnd 7.200510904745402u
r285 n181 Vsource 2.399251954308758
c285 Vsource gnd 7.200510904745402u
r289 n157 Vsource 2.399251954308758
c289 Vsource gnd 7.200510904745402u
r291 n175 Vsource 2.399251954308758
c291 Vsource gnd 7.200510904745402u
r295 n146 Vsource 2.399251954308758
c295 Vsource gnd 7.200510904745402u
r296 n140 Vsource 2.399251954308758
c296 Vsource gnd 7.200510904745402u
r297 n129 Vsource 2.399251954308758
c297 Vsource gnd 7.200510904745402u
r298 n120 Vsource 2.399251954308758
c298 Vsource gnd 7.200510904745402u
r299 n200 Vsource 2.399251954308758
c299 Vsource gnd 7.200510904745402u
r300 n144 Vsource 2.399251954308758
c300 Vsource gnd 7.200510904745402u
r301 n187 Vsource 2.399251954308758
c301 Vsource gnd 7.200510904745402u
r302 n122 Vsource 2.399251954308758
c302 Vsource gnd 7.200510904745402u
r304 n144 Vsource 2.399251954308758
c304 Vsource gnd 7.200510904745402u
r305 n172 Vsource 2.399251954308758
c305 Vsource gnd 7.200510904745402u
r307 n117 Vsource 2.399251954308758
c307 Vsource gnd 7.200510904745402u
r309 n141 Vsource 2.399251954308758
c309 Vsource gnd 7.200510904745402u
r311 n161 Vsource 2.399251954308758
c311 Vsource gnd 7.200510904745402u
r312 n152 Vsource 2.399251954308758
c312 Vsource gnd 7.200510904745402u
r313 n199 Vsource 2.399251954308758
c313 Vsource gnd 7.200510904745402u
r315 n139 Vsource 2.399251954308758
c315 Vsource gnd 7.200510904745402u
r317 n194 Vsource 2.399251954308758
c317 Vsource gnd 7.200510904745402u
r319 n188 Vsource 2.399251954308758
c319 Vsource gnd 7.200510904745402u
r322 n169 Vsource 2.399251954308758
c322 Vsource gnd 7.200510904745402u
r323 n130 Vsource 2.399251954308758
c323 Vsource gnd 7.200510904745402u
r325 n153 Vsource 2.399251954308758
c325 Vsource gnd 7.200510904745402u
r326 n146 Vsource 2.399251954308758
c326 Vsource gnd 7.200510904745402u
r327 n155 Vsource 2.399251954308758
c327 Vsource gnd 7.200510904745402u
r330 n157 Vsource 2.399251954308758
c330 Vsource gnd 7.200510904745402u
r331 n133 Vsource 2.399251954308758
c331 Vsource gnd 7.200510904745402u
r332 n132 Vsource 2.399251954308758
c332 Vsource gnd 7.200510904745402u
r333 n142 Vsource 2.399251954308758
c333 Vsource gnd 7.200510904745402u

.end
